magic
tech scmos
magscale 1 4
timestamp 1511266102
<< metal1 >>
rect 6185 23023 6191 24023
rect 7985 23245 7991 24023
rect 9785 23467 9791 24023
rect 11585 23689 11591 24023
rect 16985 23689 16991 24023
rect 11585 23683 14669 23689
rect 9785 23461 14434 23467
rect 7985 23239 14199 23245
rect 6185 23017 13965 23023
rect 13959 15757 13965 23017
rect 14193 15757 14199 23239
rect 14428 15757 14434 23461
rect 14663 15757 14669 23683
rect 15367 23683 16991 23689
rect 15367 15757 15373 23683
rect 18785 23467 18791 24023
rect 15601 23461 18791 23467
rect 15601 15757 15607 23461
rect 20585 23245 20591 24023
rect 15836 23239 20591 23245
rect 15836 15757 15842 23239
rect 22385 23023 22391 24023
rect 16071 23017 22391 23023
rect 16071 15757 16077 23017
rect 23015 16967 24021 16973
rect 23015 15723 23021 16967
rect 16111 15717 23021 15723
rect 6142 14928 13925 14934
rect 6142 13073 6148 14928
rect 6015 13067 6148 13073
rect 13959 7023 13965 14283
rect 6165 7017 13965 7023
rect 6165 6017 6171 7017
rect 14193 6801 14199 14283
rect 7965 6795 14199 6801
rect 7965 6017 7971 6795
rect 14428 6578 14434 14283
rect 9765 6572 14434 6578
rect 9765 6017 9771 6572
rect 14663 6356 14669 14283
rect 11565 6350 14669 6356
rect 15367 6356 15373 14283
rect 15601 6578 15607 14283
rect 15836 6801 15842 14283
rect 16071 7023 16077 14283
rect 16071 7017 22371 7023
rect 15836 6795 20571 6801
rect 15601 6572 18771 6578
rect 15367 6350 16971 6356
rect 11565 6017 11571 6350
rect 16965 6017 16971 6350
rect 18765 6017 18771 6572
rect 20565 6017 20571 6795
rect 22365 6017 22371 7017
<< m2contact >>
rect 14988 16116 15004 16132
rect 15222 15952 15238 15968
rect 13550 15712 13566 15728
rect 13714 15406 13730 15422
rect 16470 15195 16486 15211
rect 16306 14312 16322 14328
rect 13786 14156 13802 14160
rect 13782 14152 13802 14156
rect 13778 14148 13802 14152
rect 13774 14144 13802 14148
rect 13770 14140 13798 14144
rect 13766 14136 13794 14140
rect 13762 14132 13790 14136
rect 13758 14128 13786 14132
rect 13754 14124 13782 14128
rect 13750 14120 13778 14124
rect 13746 14116 13774 14120
rect 13742 14112 13770 14116
rect 13738 14108 13766 14112
rect 13734 14104 13762 14108
rect 13730 14100 13758 14104
rect 13726 14096 13754 14100
rect 13722 14092 13750 14096
rect 13718 14088 13746 14092
rect 13714 14084 13742 14088
rect 13714 14080 13738 14084
rect 13714 14076 13734 14080
rect 13714 14072 13730 14076
rect 13622 13992 13638 13996
rect 13618 13988 13638 13992
rect 13614 13984 13638 13988
rect 13610 13980 13638 13984
rect 13606 13976 13634 13980
rect 13602 13972 13630 13976
rect 13598 13968 13626 13972
rect 13594 13964 13622 13968
rect 13590 13960 13618 13964
rect 13586 13956 13614 13960
rect 13582 13952 13610 13956
rect 13578 13948 13606 13952
rect 13574 13944 13602 13948
rect 13570 13940 13598 13944
rect 13566 13936 13594 13940
rect 13562 13932 13590 13936
rect 13558 13928 13586 13932
rect 13554 13924 13582 13928
rect 13550 13920 13578 13924
rect 13550 13916 13574 13920
rect 13550 13912 13570 13916
rect 13550 13908 13566 13912
<< metal2 >>
rect 7015 14317 13925 14323
rect 7015 9473 7021 14317
rect 6015 9467 7021 9473
<< metal3 >>
rect 15911 23830 15917 24031
rect 15227 23824 15917 23830
rect 14986 16114 15006 16134
rect 15227 15970 15233 23824
rect 15220 15963 15240 15970
rect 6007 15913 6575 15919
rect 6569 15417 6575 15913
rect 13719 15885 16317 15963
rect 13719 15417 13797 15885
rect 13952 15750 13972 15770
rect 14187 15750 14207 15770
rect 14421 15750 14441 15770
rect 14656 15750 14676 15770
rect 15360 15750 15380 15770
rect 15595 15750 15615 15770
rect 15829 15750 15849 15770
rect 16064 15750 16084 15770
rect 16104 15710 16124 15730
rect 6569 15411 13797 15417
rect 13719 14155 13797 15411
rect 13912 14921 13932 14941
rect 13912 14310 13932 14330
rect 16239 14323 16317 15885
rect 16239 14317 23029 14323
rect 13952 14270 13972 14290
rect 14187 14270 14207 14290
rect 14421 14270 14441 14290
rect 14656 14270 14676 14290
rect 15360 14270 15380 14290
rect 15595 14270 15615 14290
rect 15829 14270 15849 14290
rect 16064 14270 16084 14290
rect 16239 14155 16317 14317
rect 13719 14077 16317 14155
rect 23023 14127 23029 14317
rect 23023 14121 24029 14127
rect 14996 6033 15002 14077
rect 14119 6027 15002 6033
rect 14119 6009 14125 6027
<< metal4 >>
rect 14115 24010 14121 24031
rect 14115 24004 14999 24010
rect 6007 17717 7013 17723
rect 7007 15723 7013 17717
rect 14993 16127 14999 24004
rect 13555 16049 16481 16127
rect 13555 15723 13633 16049
rect 7007 15717 13633 15723
rect 13555 13991 13633 15717
rect 16403 15206 16481 16049
rect 23761 15917 24029 15923
rect 23761 15206 23767 15917
rect 16403 15200 23767 15206
rect 16403 13991 16481 15200
rect 13555 13913 16481 13991
rect 15230 6218 15236 13913
rect 15230 6212 15921 6218
rect 15915 6009 15921 6212
use PADFC  PADFC_1
timestamp 1511266102
transform 1 0 18 0 1 24020
box 0 0 6000 6000
use PADOUT  PADOUT_1
timestamp 1511266102
transform 1 0 6018 0 1 24020
box 0 0 1800 6000
use PADOUT  PADOUT_3
timestamp 1511266102
transform 1 0 7818 0 1 24020
box 0 0 1800 6000
use PADOUT  PADOUT_4
timestamp 1511266102
transform 1 0 9618 0 1 24020
box 0 0 1800 6000
use PADOUT  PADOUT_5
timestamp 1511266102
transform 1 0 11418 0 1 24020
box 0 0 1800 6000
use PADVDD  PADVDD_4
timestamp 1511266102
transform 1 0 13218 0 1 24020
box 0 0 1800 6000
use PADGND  PADGND_4
timestamp 1511266102
transform 1 0 15018 0 1 24020
box 0 0 1800 6000
use PADOUT  PADOUT_6
timestamp 1511266102
transform 1 0 16818 0 1 24020
box 0 0 1800 6000
use PADOUT  PADOUT_7
timestamp 1511266102
transform 1 0 18618 0 1 24020
box 0 0 1800 6000
use PADOUT  PADOUT_8
timestamp 1511266102
transform 1 0 20418 0 1 24020
box 0 0 1800 6000
use PADOUT  PADOUT_2
timestamp 1511266102
transform 1 0 22218 0 1 24020
box 0 0 1800 6000
use PADFC  PADFC_3
timestamp 1511266102
transform 0 1 24018 -1 0 30020
box 0 0 6000 6000
use PADNC  PADNC_2
timestamp 1511266102
transform 0 -1 6018 1 0 22220
box 0 0 1800 6000
use PADNC  PADNC_6
timestamp 1511266102
transform 0 -1 6018 1 0 20420
box 0 0 1800 6000
use PADNC  PADNC_5
timestamp 1511266102
transform 0 -1 6018 1 0 18620
box 0 0 1800 6000
use PADVDD  PADVDD_2
timestamp 1511266102
transform 0 -1 6018 1 0 16820
box 0 0 1800 6000
use PADGND  PADGND_2
timestamp 1511266102
transform 0 -1 6018 1 0 15020
box 0 0 1800 6000
use PADNC  PADNC_8
timestamp 1511266102
transform 0 1 24018 -1 0 24020
box 0 0 1800 6000
use PADNC  PADNC_13
timestamp 1511266102
transform 0 1 24018 -1 0 22220
box 0 0 1800 6000
use PADNC  PADNC_12
timestamp 1511266102
transform 0 1 24018 -1 0 20420
box 0 0 1800 6000
use PADINC  PADINC_11
timestamp 1511266102
transform 0 1 24018 -1 0 18620
box 0 0 1800 6000
use DFFPOSX1  DFFPOSX1_10
timestamp 1511266102
transform 1 0 13962 0 1 15520
box 0 0 192 200
use OAI21X1  OAI21X1_15
timestamp 1511266102
transform 1 0 14154 0 1 15520
box 0 0 64 200
use OAI21X1  OAI21X1_14
timestamp 1511266102
transform -1 0 14282 0 1 15520
box 0 0 64 200
use OAI21X1  OAI21X1_17
timestamp 1511266102
transform -1 0 14346 0 1 15520
box 0 0 64 200
use INVX1  INVX1_8
timestamp 1511266102
transform -1 0 14378 0 1 15520
box 0 0 32 200
use NOR2X1  NOR2X1_4
timestamp 1511266102
transform 1 0 14378 0 1 15520
box 0 0 48 200
use NAND2X1  NAND2X1_11
timestamp 1511266102
transform 1 0 14426 0 1 15520
box 0 0 48 200
use OAI21X1  OAI21X1_19
timestamp 1511266102
transform 1 0 14474 0 1 15520
box 0 0 64 200
use INVX1  INVX1_10
timestamp 1511266102
transform 1 0 14538 0 1 15520
box 0 0 32 200
use NOR2X1  NOR2X1_5
timestamp 1511266102
transform -1 0 14618 0 1 15520
box 0 0 48 200
use XNOR2X1  XNOR2X1_2
timestamp 1511266102
transform -1 0 14730 0 1 15520
box 0 0 112 200
use BUFX2  BUFX2_2
timestamp 1511266102
transform -1 0 14778 0 1 15520
box 0 0 48 200
use NAND2X1  NAND2X1_10
timestamp 1511266102
transform -1 0 14826 0 1 15520
box 0 0 48 200
use OAI21X1  OAI21X1_18
timestamp 1511266102
transform 1 0 14826 0 1 15520
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_2
timestamp 1511266102
transform -1 0 15082 0 1 15520
box 0 0 192 200
use DFFPOSX1  DFFPOSX1_5
timestamp 1511266102
transform 1 0 15082 0 1 15520
box 0 0 192 200
use BUFX2  BUFX2_5
timestamp 1511266102
transform 1 0 15274 0 1 15520
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_11
timestamp 1511266102
transform 1 0 15322 0 1 15520
box 0 0 192 200
use MUX2X1  MUX2X1_3
timestamp 1511266102
transform -1 0 15610 0 1 15520
box 0 0 96 200
use INVX1  INVX1_13
timestamp 1511266102
transform -1 0 15642 0 1 15520
box 0 0 32 200
use XOR2X1  XOR2X1_4
timestamp 1511266102
transform 1 0 15642 0 1 15520
box 0 0 112 200
use INVX1  INVX1_11
timestamp 1511266102
transform 1 0 15754 0 1 15520
box 0 0 32 200
use NOR2X1  NOR2X1_6
timestamp 1511266102
transform -1 0 15834 0 1 15520
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_3
timestamp 1511266102
transform 1 0 15834 0 1 15520
box 0 0 192 200
use BUFX2  BUFX2_3
timestamp 1511266102
transform 1 0 16026 0 1 15520
box 0 0 48 200
use BUFX2  BUFX2_1
timestamp 1511266102
transform -1 0 14010 0 -1 15320
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_1
timestamp 1511266102
transform -1 0 14202 0 -1 15320
box 0 0 192 200
use AND2X2  AND2X2_3
timestamp 1511266102
transform -1 0 14266 0 -1 15320
box 0 0 64 200
use INVX1  INVX1_6
timestamp 1511266102
transform 1 0 14266 0 -1 15320
box 0 0 32 200
use OAI21X1  OAI21X1_16
timestamp 1511266102
transform -1 0 14362 0 -1 15320
box 0 0 64 200
use NAND2X1  NAND2X1_9
timestamp 1511266102
transform -1 0 14410 0 -1 15320
box 0 0 48 200
use INVX1  INVX1_5
timestamp 1511266102
transform -1 0 14442 0 -1 15320
box 0 0 32 200
use DFFPOSX1  DFFPOSX1_9
timestamp 1511266102
transform -1 0 14634 0 -1 15320
box 0 0 192 200
use MUX2X1  MUX2X1_4
timestamp 1511266102
transform 1 0 14634 0 -1 15320
box 0 0 96 200
use DFFPOSX1  DFFPOSX1_13
timestamp 1511266102
transform 1 0 14730 0 -1 15320
box 0 0 192 200
use MUX2X1  MUX2X1_2
timestamp 1511266102
transform -1 0 15018 0 -1 15320
box 0 0 96 200
use INVX1  INVX1_3
timestamp 1511266102
transform -1 0 15050 0 -1 15320
box 0 0 32 200
use NOR2X1  NOR2X1_1
timestamp 1511266102
transform 1 0 15050 0 -1 15320
box 0 0 48 200
use OAI22X1  OAI22X1_1
timestamp 1511266102
transform 1 0 15098 0 -1 15320
box 0 0 80 200
use INVX1  INVX1_1
timestamp 1511266102
transform -1 0 15210 0 -1 15320
box 0 0 32 200
use XOR2X1  XOR2X1_1
timestamp 1511266102
transform 1 0 15210 0 -1 15320
box 0 0 112 200
use OAI21X1  OAI21X1_2
timestamp 1511266102
transform -1 0 15386 0 -1 15320
box 0 0 64 200
use OAI21X1  OAI21X1_20
timestamp 1511266102
transform -1 0 15450 0 -1 15320
box 0 0 64 200
use NAND2X1  NAND2X1_12
timestamp 1511266102
transform 1 0 15450 0 -1 15320
box 0 0 48 200
use NAND3X1  NAND3X1_2
timestamp 1511266102
transform -1 0 15562 0 -1 15320
box 0 0 64 200
use INVX1  INVX1_12
timestamp 1511266102
transform 1 0 15562 0 -1 15320
box 0 0 32 200
use OAI22X1  OAI22X1_3
timestamp 1511266102
transform -1 0 15674 0 -1 15320
box 0 0 80 200
use OAI21X1  OAI21X1_21
timestamp 1511266102
transform -1 0 15738 0 -1 15320
box 0 0 64 200
use NOR2X1  NOR2X1_7
timestamp 1511266102
transform 1 0 15738 0 -1 15320
box 0 0 48 200
use OAI21X1  OAI21X1_1
timestamp 1511266102
transform 1 0 15786 0 -1 15320
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_4
timestamp 1511266102
transform 1 0 15850 0 -1 15320
box 0 0 192 200
use PADNC  PADNC_4
timestamp 1511266102
transform 0 -1 6018 1 0 13220
box 0 0 1800 6000
use PADVDD  PADVDD_3
timestamp 1511266102
transform 0 1 24018 -1 0 16820
box 0 0 1800 6000
use DFFPOSX1  DFFPOSX1_14
timestamp 1511266102
transform 1 0 13962 0 1 14720
box 0 0 192 200
use OAI21X1  OAI21X1_11
timestamp 1511266102
transform 1 0 14154 0 1 14720
box 0 0 64 200
use OAI21X1  OAI21X1_10
timestamp 1511266102
transform -1 0 14282 0 1 14720
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_15
timestamp 1511266102
transform 1 0 14282 0 1 14720
box 0 0 192 200
use MUX2X1  MUX2X1_1
timestamp 1511266102
transform -1 0 14570 0 1 14720
box 0 0 96 200
use BUFX2  BUFX2_6
timestamp 1511266102
transform -1 0 14618 0 1 14720
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_6
timestamp 1511266102
transform -1 0 14810 0 1 14720
box 0 0 192 200
use XOR2X1  XOR2X1_2
timestamp 1511266102
transform 1 0 14810 0 1 14720
box 0 0 112 200
use INVX1  INVX1_4
timestamp 1511266102
transform 1 0 14922 0 1 14720
box 0 0 32 200
use INVX1  INVX1_2
timestamp 1511266102
transform 1 0 14954 0 1 14720
box 0 0 32 200
use OAI21X1  OAI21X1_4
timestamp 1511266102
transform 1 0 14986 0 1 14720
box 0 0 64 200
use NAND2X1  NAND2X1_4
timestamp 1511266102
transform -1 0 15098 0 1 14720
box 0 0 48 200
use OAI22X1  OAI22X1_2
timestamp 1511266102
transform 1 0 15098 0 1 14720
box 0 0 80 200
use AOI21X1  AOI21X1_3
timestamp 1511266102
transform 1 0 15178 0 1 14720
box 0 0 64 200
use OAI21X1  OAI21X1_3
timestamp 1511266102
transform -1 0 15306 0 1 14720
box 0 0 64 200
use OR2X2  OR2X2_1
timestamp 1511266102
transform -1 0 15370 0 1 14720
box 0 0 64 200
use AND2X2  AND2X2_2
timestamp 1511266102
transform -1 0 15434 0 1 14720
box 0 0 64 200
use NAND2X1  NAND2X1_2
timestamp 1511266102
transform 1 0 15434 0 1 14720
box 0 0 48 200
use AOI21X1  AOI21X1_2
timestamp 1511266102
transform -1 0 15546 0 1 14720
box 0 0 64 200
use NAND2X1  NAND2X1_1
timestamp 1511266102
transform -1 0 15594 0 1 14720
box 0 0 48 200
use INVX1  INVX1_9
timestamp 1511266102
transform 1 0 15594 0 1 14720
box 0 0 32 200
use NOR2X1  NOR2X1_3
timestamp 1511266102
transform -1 0 15674 0 1 14720
box 0 0 48 200
use INVX1  INVX1_7
timestamp 1511266102
transform -1 0 15706 0 1 14720
box 0 0 32 200
use NAND2X1  NAND2X1_14
timestamp 1511266102
transform 1 0 15706 0 1 14720
box 0 0 48 200
use AOI21X1  AOI21X1_5
timestamp 1511266102
transform -1 0 15818 0 1 14720
box 0 0 64 200
use AOI21X1  AOI21X1_1
timestamp 1511266102
transform 1 0 15818 0 1 14720
box 0 0 64 200
use AND2X2  AND2X2_1
timestamp 1511266102
transform -1 0 15946 0 1 14720
box 0 0 64 200
use XOR2X1  XOR2X1_5
timestamp 1511266102
transform 1 0 15946 0 1 14720
box 0 0 112 200
use DFFPOSX1  DFFPOSX1_16
timestamp 1511266102
transform 1 0 13962 0 -1 14520
box 0 0 192 200
use OAI21X1  OAI21X1_9
timestamp 1511266102
transform 1 0 14154 0 -1 14520
box 0 0 64 200
use OAI21X1  OAI21X1_8
timestamp 1511266102
transform -1 0 14282 0 -1 14520
box 0 0 64 200
use BUFX2  BUFX2_7
timestamp 1511266102
transform -1 0 14330 0 -1 14520
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_7
timestamp 1511266102
transform -1 0 14522 0 -1 14520
box 0 0 192 200
use XOR2X1  XOR2X1_3
timestamp 1511266102
transform 1 0 14522 0 -1 14520
box 0 0 112 200
use NAND2X1  NAND2X1_7
timestamp 1511266102
transform 1 0 14634 0 -1 14520
box 0 0 48 200
use NAND2X1  NAND2X1_3
timestamp 1511266102
transform 1 0 14682 0 -1 14520
box 0 0 48 200
use OAI21X1  OAI21X1_6
timestamp 1511266102
transform -1 0 14794 0 -1 14520
box 0 0 64 200
use NOR2X1  NOR2X1_2
timestamp 1511266102
transform 1 0 14794 0 -1 14520
box 0 0 48 200
use OR2X2  OR2X2_2
timestamp 1511266102
transform -1 0 14906 0 -1 14520
box 0 0 64 200
use OAI21X1  OAI21X1_5
timestamp 1511266102
transform -1 0 14970 0 -1 14520
box 0 0 64 200
use NAND2X1  NAND2X1_5
timestamp 1511266102
transform -1 0 15018 0 -1 14520
box 0 0 48 200
use XNOR2X1  XNOR2X1_1
timestamp 1511266102
transform 1 0 15018 0 -1 14520
box 0 0 112 200
use NAND3X1  NAND3X1_1
timestamp 1511266102
transform -1 0 15194 0 -1 14520
box 0 0 64 200
use AOI21X1  AOI21X1_4
timestamp 1511266102
transform 1 0 15194 0 -1 14520
box 0 0 64 200
use NAND2X1  NAND2X1_8
timestamp 1511266102
transform -1 0 15306 0 -1 14520
box 0 0 48 200
use OAI21X1  OAI21X1_7
timestamp 1511266102
transform 1 0 15306 0 -1 14520
box 0 0 64 200
use NAND2X1  NAND2X1_6
timestamp 1511266102
transform -1 0 15418 0 -1 14520
box 0 0 48 200
use BUFX2  BUFX2_8
timestamp 1511266102
transform 1 0 15418 0 -1 14520
box 0 0 48 200
use DFFPOSX1  DFFPOSX1_8
timestamp 1511266102
transform -1 0 15658 0 -1 14520
box 0 0 192 200
use OAI21X1  OAI21X1_12
timestamp 1511266102
transform 1 0 15658 0 -1 14520
box 0 0 64 200
use OAI21X1  OAI21X1_13
timestamp 1511266102
transform -1 0 15786 0 -1 14520
box 0 0 64 200
use DFFPOSX1  DFFPOSX1_12
timestamp 1511266102
transform 1 0 15786 0 -1 14520
box 0 0 192 200
use NAND2X1  NAND2X1_13
timestamp 1511266102
transform -1 0 16026 0 -1 14520
box 0 0 48 200
use BUFX2  BUFX2_4
timestamp 1511266102
transform 1 0 16026 0 -1 14520
box 0 0 48 200
use PADINC  PADINC_10
timestamp 1511266102
transform 0 -1 6018 1 0 11420
box 0 0 1800 6000
use PADNC  PADNC_3
timestamp 1511266102
transform 0 -1 6018 1 0 9620
box 0 0 1800 6000
use PADINC  PADINC_9
timestamp 1511266102
transform 0 -1 6018 1 0 7820
box 0 0 1800 6000
use PADNC  PADNC_1
timestamp 1511266102
transform 0 -1 6018 1 0 6020
box 0 0 1800 6000
use PADGND  PADGND_3
timestamp 1511266102
transform 0 1 24018 -1 0 15020
box 0 0 1800 6000
use PADNC  PADNC_11
timestamp 1511266102
transform 0 1 24018 -1 0 13220
box 0 0 1800 6000
use PADNC  PADNC_10
timestamp 1511266102
transform 0 1 24018 -1 0 11420
box 0 0 1800 6000
use PADNC  PADNC_9
timestamp 1511266102
transform 0 1 24018 -1 0 9620
box 0 0 1800 6000
use PADNC  PADNC_7
timestamp 1511266102
transform 0 1 24018 -1 0 7820
box 0 0 1800 6000
use PADFC  PADFC_2
timestamp 1511266102
transform 0 -1 6018 1 0 20
box 0 0 6000 6000
use PADINC  PADINC_1
timestamp 1511266102
transform -1 0 7818 0 -1 6020
box 0 0 1800 6000
use PADINC  PADINC_3
timestamp 1511266102
transform -1 0 9618 0 -1 6020
box 0 0 1800 6000
use PADINC  PADINC_4
timestamp 1511266102
transform -1 0 11418 0 -1 6020
box 0 0 1800 6000
use PADINC  PADINC_5
timestamp 1511266102
transform -1 0 13218 0 -1 6020
box 0 0 1800 6000
use PADGND  PADGND_1
timestamp 1511266102
transform -1 0 15018 0 -1 6020
box 0 0 1800 6000
use PADVDD  PADVDD_1
timestamp 1511266102
transform -1 0 16818 0 -1 6020
box 0 0 1800 6000
use PADINC  PADINC_6
timestamp 1511266102
transform -1 0 18618 0 -1 6020
box 0 0 1800 6000
use PADINC  PADINC_7
timestamp 1511266102
transform -1 0 20418 0 -1 6020
box 0 0 1800 6000
use PADINC  PADINC_8
timestamp 1511266102
transform -1 0 22218 0 -1 6020
box 0 0 1800 6000
use PADINC  PADINC_2
timestamp 1511266102
transform -1 0 24018 0 -1 6020
box 0 0 1800 6000
use PADFC  PADFC_4
timestamp 1511266102
transform -1 0 30018 0 -1 6020
box 0 0 6000 6000
<< labels >>
flabel metal3 14421 15750 14441 15770 6 FreeSans 48 0 0 0 q<2>
port 0 nsew
flabel metal3 14656 15750 14676 15770 6 FreeSans 48 0 0 0 q<3>
port 1 nsew
flabel metal3 16104 15710 16124 15730 6 FreeSans 48 0 0 0 e
port 2 nsew
flabel metal3 15360 14270 15380 14290 6 FreeSans 48 0 0 0 d<4>
port 3 nsew
flabel metal3 13912 14310 13932 14330 6 FreeSans 48 0 0 0 clk
port 4 nsew
flabel metal3 15829 14270 15849 14290 6 FreeSans 48 0 0 0 d<6>
port 5 nsew
flabel metal3 15829 15750 15849 15770 6 FreeSans 48 0 0 0 q<6>
port 6 nsew
flabel metal3 13952 15750 13972 15770 6 FreeSans 48 0 0 0 q<0>
port 7 nsew
flabel metal3 14187 15750 14207 15770 6 FreeSans 48 0 0 0 q<1>
port 8 nsew
flabel metal3 16064 14270 16084 14290 6 FreeSans 48 0 0 0 d<7>
port 9 nsew
flabel metal3 15360 15750 15380 15770 6 FreeSans 48 0 0 0 q<4>
port 10 nsew
flabel metal3 15595 15750 15615 15770 6 FreeSans 48 0 0 0 q<5>
port 11 nsew
flabel metal3 14656 14270 14676 14290 6 FreeSans 48 0 0 0 d<3>
port 12 nsew
flabel metal3 16064 15750 16084 15770 6 FreeSans 48 0 0 0 q<7>
port 13 nsew
flabel metal3 14986 16114 15006 16134 6 FreeSans 48 0 0 0 vdd
port 14 nsew
flabel metal3 15220 15950 15240 15970 6 FreeSans 48 0 0 0 gnd
port 15 nsew
flabel metal3 14187 14270 14207 14290 6 FreeSans 48 0 0 0 d<1>
port 16 nsew
flabel metal3 13952 14270 13972 14290 6 FreeSans 48 0 0 0 d<0>
port 17 nsew
flabel metal3 14421 14270 14441 14290 6 FreeSans 48 0 0 0 d<2>
port 18 nsew
flabel metal3 13912 14921 13932 14941 6 FreeSans 48 0 0 0 clr
port 19 nsew
flabel metal3 15595 14270 15615 14290 6 FreeSans 48 0 0 0 d<5>
port 20 nsew
<< end >>
